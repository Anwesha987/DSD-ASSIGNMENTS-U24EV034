module full_adder_tb;

    // Inputs
    reg a;
    reg b;
    reg cin;

    // Outputs
    wire sum;
    wire cout;

    // Instantiate the full adder
    full_adder uut (
        .a(a),
        .b(b),
        .cin(cin),
        .sum(sum),
        .cout(cout)
    );

  	 initial begin
        $dumpfile("output.vcd");
        $dumpvars;
     end

    // Test all combinations
    initial begin
        $display("A B Cin | Sum Cout");
        $display("--------|----------");
        a = 0; b = 0; cin = 0; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 0; b = 0; cin = 1; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 0; b = 1; cin = 0; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 0; b = 1; cin = 1; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 1; b = 0; cin = 0; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 1; b = 0; cin = 1; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 1; b = 1; cin = 0; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        a = 1; b = 1; cin = 1; #10; $display("%b %b  %b  |  %b    %b", a, b, cin, sum, cout);
        $finish;
    end

endmodule
